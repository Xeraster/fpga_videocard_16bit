`include "fifo_bram.v"
`include "managedVramDataBuffer.v"

`default_nettype none

//generate a 640x480 vga sync signal
module generateSync(
    input clock,
    output reg HSYNC,
    output reg VSYNC,
    output reg [19:0] vramAddress,
    input RESET,                 //gotta tell those counters when to reset to zero
    output reg VALID_PIXELS,             //its a 1 if there is allowed to be data on R,G,B
    output reg[10:0] horizontalCount,
    output reg[9:0] verticalCount 
);
    //reg [10:0] horizontalCount;
    //reg [9:0] verticalCount;
    reg VALID_H;                    //1 if in valid horizontal viewing area. 0 if otherwise 
    reg VALID_V;                    //1 if in valid veritcal viewing area. 0 if otherwise
    always@(posedge clock or negedge RESET)
    begin
        if (!RESET)
        begin
            horizontalCount <= 0;
            verticalCount <= 0;
            vramAddress <= 0;
        end
        else begin
        //increment h counter
        horizontalCount <= horizontalCount + 1;

        //horizontal counter cases
        if (horizontalCount >= 640 & horizontalCount < 656)
            begin
                //front porch
                VALID_H <= 0;
                HSYNC <= 1;
            end
        else if (horizontalCount >= 656 & horizontalCount < 752)
            begin
                //when hsync happens
                VALID_H <= 0;
                HSYNC <= 0;
            end
        else if (horizontalCount >= 752 & horizontalCount < 799)
            begin
                //back porch
                HSYNC <= 1;
                VALID_H <= 0;
            end
        else if (horizontalCount >= 799)
            begin
                //the reset pixel
                verticalCount <= verticalCount + 1;
                horizontalCount <= 0;
                HSYNC <= 1;
                VALID_H <= 1;
            end
        else
            begin
                //this should only be happening if within visible screen area
                HSYNC <= 1;
                VALID_H <= 1;
                vramAddress <= vramAddress + 2;
            end

        if (verticalCount >= 480 & verticalCount < 490)
            begin
                //front porch
                VALID_V <= 0;
                VSYNC <= 1;
            end
        else if (verticalCount >= 490 & verticalCount < 492)
            begin
                //vsync signal
                VALID_V <= 0;
                VSYNC <= 0;
            end
        else if (verticalCount >= 492 & verticalCount < 525)
            begin
                //back porch
                VALID_V <= 0;
                VSYNC <= 1;
            end
        else if (verticalCount >= 525)
            begin
                //the reset pixel
                VALID_V <= 0;
                VSYNC <= 1;
                verticalCount <= 0;
                vramAddress <= 0;
            end
        else
            begin
                //this should only be happening if within visible screen area
                VALID_V <= 1;
                VSYNC <= 1;
            end

        //set the value of the valid pixel signal. only draw pixels if h and v are within a valid range
        VALID_PIXELS <= VALID_H & VALID_V;
        end

    end

endmodule

module tb();
reg clk;
reg rst_n;

//reg[15:0] dataIn;
wire read_en;
wire write_en;
wire[15:0] dataOut;  //wire on hardware, reg for testbench because thats just how
wire full, empty, valid;
reg[15:0] vramDataBus;
wire[15:0] vgaDataPixel;
wire[19:0] genVramAddress;       //what vram address to request
wire[19:0] maxVramAddress;
wire WE, CE, RD, done;
reg vblank;
reg pixelClock;
wire HSYNC, VSYNC, VALID_PIXELS;
wire[10:0] horizontalCount;
wire[9:0] verticalCount;
wire[19:0] vramAddress;

reg bus_free;

wire[4:0] Ri;
wire[5:0] Gi;
wire[4:0] Bi;
wire frameEnd;
wire almostFull;

assign maxVramAddress = 20'h96000;

localparam PIXELCLK_PERIOD = 10;
localparam CLK_PERIOD = 4;
always #(CLK_PERIOD/2) clk=~clk;

generateSync gsc(pixelClock, HSYNC, VSYNC, vramAddress, rst_n, VALID_PIXELS, horizontalCount, verticalCount);

//bram_256x16 testram(dataIn, write_en, waddr, clk, raddr, clk, dataOut);
psuedofiforam testfifo(vramDataBus, write_en, read_en, ~clk, pixelClock, dataOut, rst_n, full, empty, valid, almostFull);
managedVramDataBuffer testramthingy(vramDataBus, Ri, Gi, Bi, RD, CE, clk, done, bus_free, VALID_PIXELS, empty, full, valid, write_en, read_en, genVramAddress, maxVramAddress, rst_n, pixelClock, dataOut, frameEnd, almostFull);

initial begin
    $dumpfile("tb_.vcd");
    $dumpvars(0, tb); 
end

initial begin
    #1 rst_n<=1'bx;clk<=1'bx;
    #(CLK_PERIOD*3) rst_n<=1;
    #(CLK_PERIOD*3) rst_n<=0;clk<=0;
    repeat(20) @(posedge clk);
    rst_n<=1;
    @(posedge clk);
    repeat(10000) @(posedge clk);
    $finish(2);
end

initial begin
    #(PIXELCLK_PERIOD)
    bus_free = 0;
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    bus_free = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    bus_free=0;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
    #(PIXELCLK_PERIOD)
    pixelClock = 1;
    #(PIXELCLK_PERIOD)
    pixelClock = 0;
end

initial begin
    //ugh
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
    #(CLK_PERIOD)
    vramDataBus=420;
    #(CLK_PERIOD)
    vramDataBus=4442;
    #(CLK_PERIOD)
    vramDataBus=55555;
    #(CLK_PERIOD)
    vramDataBus=1234;
    #(CLK_PERIOD)
    vramDataBus=69;
    #(CLK_PERIOD)
    vramDataBus=6996;
end

endmodule
