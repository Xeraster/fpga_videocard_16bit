`include "writeBufferVram_different.v"

`default_nettype none

module bram_256x16(din, write_en, waddr, wclk, raddr, rclk, dout);//256x16
parameter addr_width = 8;
parameter data_width = 16;
input [addr_width-1:0] waddr, raddr;
input [data_width-1:0] din;
input write_en, wclk, rclk;
output reg [data_width-1:0] dout;
reg [data_width-1:0] mem [(1<<addr_width)-1:0];

always @(posedge wclk) // Write memory.
begin
    if (write_en)
    begin
        mem[waddr] <= din; // Using write address bus.
    end
end

always @(posedge rclk) // Read memory.
begin
    dout <= mem[raddr]; // Using read address bus.
end
endmodule

module tb();
reg clk;
reg readClk;
reg rst_n;
reg test_signal;

reg[15:0] dataIn;
reg[19:0] addressFromIsa;
wire[15:0] dataOut;
wire [19:0] addressOut;
wire full, almostFull, WRITEBUF_IO_EN, empty;
wire write_cmd, chip_select;
reg bus_free;
reg newData;//on the rising edge of this, it writes to the write buffer
localparam CLK_PERIOD = 6;
localparam READCLK_PERIOD = 10;
always #(CLK_PERIOD/2) clk=~clk;

//bram_256x16 testram(dataIn, write_en, waddr, clk, raddr, clk, dataOut);
writeBufferVram testWriteBuffer(dataIn, addressFromIsa, clk, newData, dataOut, addressOut, write_cmd, chip_select, bus_free, readClk, rst_n, WRITEBUF_IO_EN, full, almostFull, empty);

initial begin
    $dumpfile("tb_.vcd");
    $dumpvars(0, tb);
end

/*initial begin
    #1 rst_n<=1'bx;clk<=1'bx;
    #(CLK_PERIOD*3) rst_n<=1;
    #(CLK_PERIOD*3) rst_n<=0;clk<=0;
    repeat(2) @(posedge clk);
    rst_n<=1;
    @(posedge clk);
    repeat(10) @(posedge clk);
    $finish(2);
end*/
//too difficult to control

initial begin
    #(CLK_PERIOD/2)
    bus_free=1;
    newData=0;
    dataIn=16'h420;
    addressFromIsa=16'h0;
    rst_n=1;
    clk=1;
    #(CLK_PERIOD/2)
    clk=0;
    #(CLK_PERIOD/2)
    clk=1;
    rst_n=0;
    #(CLK_PERIOD/2)
    clk=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=1;
    #(CLK_PERIOD/2)
    clk=1;
    rst_n=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    #(CLK_PERIOD/2)
    clk=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    newData=0;
    #(CLK_PERIOD/2)
    clk=1;
    newData=1;
    #(CLK_PERIOD/2)
    clk=0;
    #(CLK_PERIOD/2)
    clk=1;
    #(CLK_PERIOD/2)
    clk=0;
    #(CLK_PERIOD/2)
    clk=1;
    #(CLK_PERIOD/2)
    clk=0;
end

initial begin
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    #(READCLK_PERIOD/2)
    readClk=1;
    #(READCLK_PERIOD/2)
    readClk=0;
    $finish(2);
end

endmodule
